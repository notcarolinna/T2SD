module timer 
(
  // Declarar os pinos de IO
);

endmodule