module timer 
(
  input 
);

endmodule
