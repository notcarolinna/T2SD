module dcm 
(
  // Declarar os pinos I/O
);

endmodule